`timescale 1ns / 1ps

module addsub4b(add_sub, A3, A2, A1, A0, B3, B2, B1, B0, Co, R3, R2, R1, R0);
  input add_sub;  // Se add_sub=0 faz A+B; se add_sub=1 faz A-B
  input A3, A2, A1, A0;  // Operando A
  input B3, B2, B1, B0;  // Operando B 
  output Co;
  output R3, R2, R1, R0; // Resultado R

  // Acrescente a seguir a implementa��o

  
  
endmodule
